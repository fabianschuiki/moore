package foo is
	alias bar is baz;
	alias bar is baz [];
	alias bar is baz [a,b,c];
	alias bar is baz [return d];
	alias bar is baz [a,b,c return d];
end;
