entity foo is end;
architecture bar of foo is

	constant A : std.standard.BOOLEAN;
	constant B : BOOLEAN := FALSE;
	constant C : BOOLEAN := TRUE;

begin end;
