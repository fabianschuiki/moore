module A;
    for (genvar i = 0; i < 4; i++)
        B b();
endmodule

module B;
endmodule
