module mh4 (var x); // ERROR: direction defaults to inout, which cannot be var
endmodule
