entity foo is end;
architecture bar of foo is

	constant A : std.standard.BIT;
	constant B : BIT := '0';
	constant C : BIT := '1';

begin end;
