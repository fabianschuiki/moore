entity foo is end;
architecture bar of foo is

	constant xA : std.standard.TIME;
	--constant xB : TIME := 10 ns;

	--constant yA: std.standard.DELAY_LENGTH;

	--constant zA: std.standard.TIME_VECTOR;

begin end;
