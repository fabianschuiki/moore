(* dont_touch = "true" *)
