// RUN: moore %s -e foo -Vinsts

module foo;
endmodule
