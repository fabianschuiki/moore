module a0;
	logic [3:0] a;
	logic [8:0] b;

	assign a = (b + 2) - '1;
endmodule
