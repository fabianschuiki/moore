module a0;
	logic [15:0] x, y;

	initial begin
		if (x);
		while (x);
		do begin
		end while (x);
	end
endmodule
