module A;
	int a;
	initial;
	initial a = 42;
endmodule
