module a0;
	bit [15:0] x;
	bit [63:0] y;
	assign y = 32'(x);
endmodule
