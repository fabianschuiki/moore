module A;
	int a;
	initial a = 42;
endmodule
