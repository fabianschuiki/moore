// RUN: moore %s -e foo -O0

module foo;
	bar x();
	logic z;
	assign z = x.valid & x.ready | !x.data;
endmodule

interface bar;
	logic [31:0] data;
	logic valid;
	logic ready;
endinterface

// CHECK: entity @foo () -> () {
// CHECK:     %x.data = sig i32 %1
// CHECK:     %x.valid = sig i1 %2
// CHECK:     %x.ready = sig i1 %3
// CHECK:     %4 = and i1 %x.valid1, %x.ready1
// CHECK:     %6 = neq i32 %x.data1, %5
// CHECK: }
