-- This file tests sequential statements.
