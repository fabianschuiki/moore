module A;
endmodule

module B (
	input bit x,
	output bit y,
	inout bit z
);
endmodule
